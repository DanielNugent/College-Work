library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity memory is 
    Port(
        address : in std_logic_vector(15 downto 0);
        WD : in std_logic_vector(15 downto 0); --in
        MW : in std_logic;
        MR : in std_logic;
        read_data : out std_logic_vector(15 downto 0) -- out
    );
end memory;


architecture Behavioral of memory is
    type mem_array is array(0 to 511) of std_logic_vector(15 downto 0);
    -- define type, for memory arrays
begin

    mem_process : process(address, WD, MW)
    -- initialise data memory, X denotes a hexadecimal number
        variable data_mem : mem_array :=(
			x"0000", --0 
			x"0000", --1 store in reg 0
			x"0241", --2 store in reg 1
			x"0482", --3 store in reg 2
			x"06C3", --4 store in reg 3
			x"0904", --5 store in reg 4
			x"0B45", --6 store in reg 5
			x"0D86", --7 store in reg 6
			x"0FC7", --8 store in reg 7
			x"11BE", --9 ADD -> add operands
			x"1230", --A LDR -> load to r0 from memory
			x"1401", --B STR -> store from r1 into memory address
			x"1650", --C INC -> increment value in r2 by 1 and store in r1
			x"1928", --D CMP -> compliment value in r5 and store in r4
			x"1A9B", --E ADD -> adds values and stores into r2 via r3
			x"1C52", --F BCH -> branch unconditionally
			
			--module 01
			x"2652", --0 ADD STR r1 -> add and store into r1
			x"2802", --1 BCZ -> branch conditionally if z is set thereby skipping the next add instruction
			x"2A5B", --2 ADD STR r1 -> add and stores into r1
			x"2D9B", --3 ADD STR r6 -> add and stores into r6
			x"2F9B", --4 ADD STR r6 -> add and stores into r6
		
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            -- 64
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            -- 128
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            -- 192
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            -- 256
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            -- 320
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            -- 384
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            -- 448
           
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000", x"0000",
            x"0000", x"0000", x"0000"
            -- 512
        );

       	variable addr : integer range 0 to 511;
        variable addr_out : STD_LOGIC_VECTOR(15 downto 0);
        
        begin
            addr := conv_integer(address(8 downto 0));
            addr_out := data_mem(addr);
            if MW = '1' then
                data_mem(addr) := WD;
            else read_data <= addr_out;
            end if;
        end process;


end Behavioral ; -- Behavioral

